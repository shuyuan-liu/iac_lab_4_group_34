module f1_cpu #(
    parameter ADDR_WIDTH = 16,
              DATA_WIDTH = 32
)(
   input logic clk,
   output logic a0,

)
