module adder(
    input [31:0] i1,
    input [31:0] i2,
    output [31:0] out
);

assign out = i1 + i2;

endmodule
